library verilog;
use verilog.vl_types.all;
entity tb1 is
end tb1;
